
module counter(
	input logic increment, 
	input logic reset,
	input logic clk,
	output logic [3:0]
);

logic input [3:0] next_state;

always_comb
	if (increment)
		next_state = 
end


always_ff

end



endmodule
