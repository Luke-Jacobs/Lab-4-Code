
module multiplier_fsm(
	input logic reset,
	input logic clk,
	input logic run,
	input logic clearA_loadB,
	output logic shift,
	output logic add,
	output logic sub
);

always_comb

end

always_ff

end


endmodule
